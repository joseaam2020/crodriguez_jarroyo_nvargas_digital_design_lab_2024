// spi_master.v

// Generated using ACDS version 20.1 711

`timescale 1 ps / 1 ps
module spi_master (
		input  wire        spi_0_clk_clk,                     //              spi_0_clk.clk
		input  wire        spi_0_external_MISO,               //         spi_0_external.MISO
		output wire        spi_0_external_MOSI,               //                       .MOSI
		output wire        spi_0_external_SCLK,               //                       .SCLK
		output wire        spi_0_external_SS_n,               //                       .SS_n
		output wire        spi_0_irq_irq,                     //              spi_0_irq.irq
		input  wire        spi_0_reset_reset_n,               //            spi_0_reset.reset_n
		input  wire [15:0] spi_0_spi_control_port_writedata,  // spi_0_spi_control_port.writedata
		output wire [15:0] spi_0_spi_control_port_readdata,   //                       .readdata
		input  wire [2:0]  spi_0_spi_control_port_address,    //                       .address
		input  wire        spi_0_spi_control_port_read_n,     //                       .read_n
		input  wire        spi_0_spi_control_port_chipselect, //                       .chipselect
		input  wire        spi_0_spi_control_port_write_n     //                       .write_n
	);

	spi_master_spi_master spi_master (
		.clk           (spi_0_clk_clk),                     //              clk.clk
		.reset_n       (spi_0_reset_reset_n),               //            reset.reset_n
		.data_from_cpu (spi_0_spi_control_port_writedata),  // spi_control_port.writedata
		.data_to_cpu   (spi_0_spi_control_port_readdata),   //                 .readdata
		.mem_addr      (spi_0_spi_control_port_address),    //                 .address
		.read_n        (spi_0_spi_control_port_read_n),     //                 .read_n
		.spi_select    (spi_0_spi_control_port_chipselect), //                 .chipselect
		.write_n       (spi_0_spi_control_port_write_n),    //                 .write_n
		.irq           (spi_0_irq_irq),                     //              irq.irq
		.MISO          (spi_0_external_MISO),               //         external.export
		.MOSI          (spi_0_external_MOSI),               //                 .export
		.SCLK          (spi_0_external_SCLK),               //                 .export
		.SS_n          (spi_0_external_SS_n)                //                 .export
	);

endmodule
